--
-- entity name: g31_7_Segment_Decoder
--
-- Copyright (C) 2016 g31
-- Version 1.0
-- Author: Andrei Purcarus Vlastimil Lacina
-- Date: October 6th, 2016

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY g31_7_Segment_Decoder IS
	PORT (
		ASCII_CODE : IN  STD_LOGIC_VECTOR(6 DOWNTO 0);
		SEGMENTS   : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END g31_7_Segment_Decoder;

ARCHITECTURE bdf_type OF g31_7_Segment_Decoder IS
BEGIN
	WITH ASCII_CODE SELECT
		SEGMENTS <=
			"1000000" WHEN "0110000",
			"1111001" WHEN "0110001",
			"0100100" WHEN "0110010",
			"0110000" WHEN "0110011",
			"0011001" WHEN "0110100",
			"0010010" WHEN "0110101",
			"0000011" WHEN "0110110",
			"1111000" WHEN "0110111",
			"0000000" WHEN "0111000",
			"0011000" WHEN "0111001",
			
			"0001000" WHEN "1000001",
			"0000011" WHEN "1000010",
			"1000110" WHEN "1000011",
			"0100001" WHEN "1000100",
			"0000110" WHEN "1000101",
			"0001110" WHEN "1000110",
			"1000010" WHEN "1000111",
			"0001011" WHEN "1001000",
			"1111001" WHEN "1001001",
			"1100001" WHEN "1001010",
			"0001111" WHEN "1001011",
			"1000111" WHEN "1001100",
			"1001000" WHEN "1001101",
			"0101011" WHEN "1001110",
			"1000000" WHEN "1001111",
			"0001100" WHEN "1010000",
			"0100011" WHEN "1010001",
			"1001110" WHEN "1010010",
			"0010010" WHEN "1010011",
			"0000111" WHEN "1010100",
			"1000001" WHEN "1010101",
			"1011001" WHEN "1010110",
			"1100011" WHEN "1010111",
			"0001001" WHEN "1011000",
			"0010001" WHEN "1011001",
			"0100100" WHEN "1011010",
			
			"1111111" WHEN OTHERS;
END bdf_type;

