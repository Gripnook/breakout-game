--
-- entity name: g31_VGA_Test_Pattern
--
-- Copyright (C) 2016 g31
-- Version 1.0
-- Author: Andrei Purcarus Vlastimil Lacina
-- Date: October 31st, 2016

LIBRARY ieee;
USE ieee.std_logic_1164.all;
use ieee.numeric_std.all;
LIBRARY lpm;
USE lpm.lpm_components.all;

ENTITY g31_VGA_TEST_PATTERN IS
	PORT (
		CLOCK    : IN  STD_LOGIC; -- 50MHz
		RST      : IN  STD_LOGIC; -- reset
		R, G, B  : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		HSYNC    : OUT STD_LOGIC; -- horizontal sync signal
		VSYNC    : OUT STD_LOGIC -- vertical sync signal
	);
END g31_VGA_TEST_PATTERN;

ARCHITECTURE bdf_type OF g31_VGA_TEST_PATTERN IS

SIGNAL COLUMN   : UNSIGNED(9 DOWNTO 0);
SIGNAL ROW      : UNSIGNED(9 DOWNTO 0);
SIGNAL BLANKING : STD_LOGIC;

COMPONENT g31_VGA
	 PORT (
		CLOCK    : IN  STD_LOGIC; -- 50MHz
		RST      : IN  STD_LOGIC; -- reset
		BLANKING : OUT STD_LOGIC; -- blank display when zero
		ROW      : OUT UNSIGNED(9 DOWNTO 0); -- line 0 to 599
		COLUMN   : OUT UNSIGNED(9 DOWNTO 0); -- column 0 to 799
		HSYNC    : OUT STD_LOGIC; -- horizontal sync signal
		VSYNC    : OUT STD_LOGIC -- vertical sync signal
	);
END COMPONENT;

BEGIN
VGA1: g31_VGA PORT MAP (CLOCK => CLOCK, RST => RST, BLANKING => BLANKING,
								ROW => ROW, COLUMN => COLUMN, HSYNC => HSYNC, VSYNC => VSYNC);

R <=  "0000" WHEN BLANKING = '0' ELSE
		"1111" WHEN COLUMN <=  99  ELSE
		"1111" WHEN COLUMN <= 199  ELSE
		"0000" WHEN COLUMN <= 299  ELSE
		"0000" WHEN COLUMN <= 399  ELSE	
		"1111" WHEN COLUMN <= 499  ELSE
		"1111" WHEN COLUMN <= 599  ELSE
		"0000" WHEN COLUMN <= 699  ELSE
		"0000";
		
G <=  "0000" WHEN BLANKING = '0' ELSE
		"1111" WHEN COLUMN <=  99  ELSE
		"1111" WHEN COLUMN <= 199  ELSE
		"1111" WHEN COLUMN <= 299  ELSE
		"1111" WHEN COLUMN <= 399  ELSE
		"0000" WHEN COLUMN <= 499  ELSE
		"0000" WHEN COLUMN <= 599  ELSE
		"0000" WHEN COLUMN <= 699  ELSE
		"0000";
		
B <=  "0000" WHEN BLANKING = '0' ELSE
		"1111" WHEN COLUMN <=  99  ELSE
		"0000" WHEN COLUMN <= 199  ELSE
		"1111" WHEN COLUMN <= 299  ELSE
		"0000" WHEN COLUMN <= 399  ELSE
		"1111" WHEN COLUMN <= 499  ELSE
		"0000" WHEN COLUMN <= 599  ELSE
		"1111" WHEN COLUMN <= 699  ELSE
		"0000";

END bdf_type;

