--
-- entity name: g31_64_6_Encoder
--
-- Copyright (C) 2016 g31
-- Version 1.0
-- Author: Andrei Purcarus Vlastimil Lacina
-- Date: October 3rd, 2016

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY g31_64_6_Encoder IS
	PORT (
		INPUTS : IN  STD_LOGIC_VECTOR(63 DOWNTO 0);
		CODE   : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
		ERROR  : OUT STD_LOGIC
	);
END g31_64_6_Encoder;

ARCHITECTURE bdf_type OF g31_64_6_Encoder IS

COMPONENT g31_16_4_Encoder
	PORT(
		BLOCK_COL : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		CODE      : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		ERROR     : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL CODE1, CODE2, CODE3, CODE4     : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL ERROR1, ERROR2, ERROR3, ERROR4 : STD_LOGIC;

BEGIN
	ENC1 : g31_16_4_Encoder
		PORT MAP (
			BLOCK_COL => INPUTS(15 DOWNTO 0),
			CODE => CODE1,
			ERROR => ERROR1
		);
	ENC2 : g31_16_4_Encoder
		PORT MAP (
			BLOCK_COL => INPUTS(31 DOWNTO 16),
			CODE => CODE2,
			ERROR => ERROR2
		);
	ENC3 : g31_16_4_Encoder
		PORT MAP (
			BLOCK_COL => INPUTS(47 DOWNTO 32),
			CODE => CODE3,
			ERROR => ERROR3
		);
	ENC4 : g31_16_4_Encoder
		PORT MAP (
			BLOCK_COL => INPUTS(63 DOWNTO 48),
			CODE => CODE4,
			ERROR => ERROR4
		);
	CODE <=
		"000000" OR ((5 DOWNTO 4 => '0') & CODE1) WHEN ERROR1 = '0' ELSE
		"010000" OR ((5 DOWNTO 4 => '0') & CODE2) WHEN ERROR2 = '0' ELSE
		"100000" OR ((5 DOWNTO 4 => '0') & CODE3) WHEN ERROR3 = '0' ELSE
		"110000" OR ((5 DOWNTO 4 => '0') & CODE4) WHEN ERROR4 = '0' ELSE
		"000000";
	ERROR <= (ERROR1 AND ERROR2) AND (ERROR3 AND ERROR4);
END bdf_type;

